// Code your design here
class c;
  
static  reg [3:0] a;
  
  


  
endclass

module m;
  
  c c1=new();
  
  initial 
    begin 
      
      c1.a=1;
      
    end 
endmodule 
